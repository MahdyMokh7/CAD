module read_controller (
    input a, b, 
    output out
);

    assign out = a&b;

endmodule